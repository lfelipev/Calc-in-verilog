library verilog;
use verilog.vl_types.all;
entity calculadora_soma_sub_vlg_vec_tst is
end calculadora_soma_sub_vlg_vec_tst;
